----------------------------------------------------------------------------------
-- Company :         HEIA-FR
-- Engineer :        Cyril Vall�lian & Gilles Waeber
-- Module Name :     Local_display
-- Project Name :    Flappy Bird
-- Target Devices :  Spartan6
-- Description :     Local package for display constants
-- Date :            2016-06-17
-- Version :         1.0
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package local_display is
	
	type memory_m_110_30   is array(0 to 109, 0 to 29)  of std_logic_vector(7 downto 0);    -- d_score
	type memory_m_180_30   is array(0 to 179, 0 to 29)  of std_logic_vector(7 downto 0);    -- d_score_max
	type memory_m_150_30   is array(0 to 149, 0 to 29)  of std_logic_vector(7 downto 0);    -- d_title
	type memory_m_20_30    is array(0 to 19,  0 to 29)  of std_logic_vector(7 downto 0);    -- d_digit_n
	type memory_m_40_40    is array(0 to 39,  0 to 39)  of std_logic_vector(7 downto 0);    -- d_flappy
	type memory_m_40_40_bg is array(0 to 39,  0 to 39)  of std_logic;                       -- d_flappy_bg
	type memory_m_255_30   is array(0 to 254, 0 to 29)  of std_logic_vector(7 downto 0);    -- d_start_game_text
	
	
	constant d_score : memory_m_110_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"24", x"49", x"00", x"00", x"00", x"00", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"00", x"49", x"92", x"24", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"24", x"6d", x"92", x"92", x"6d", x"24", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"24", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"24", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"00", x"00", x"00", x"b6", x"92", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"00", x"00", x"00", x"b6", x"b6", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"49", x"24", x"24", x"b6", x"b6", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"24", x"24", x"24", x"24", x"b6", x"b6", x"b6", x"b6", x"24", x"24", x"24", x"24", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));

	
	constant d_score_max : memory_m_180_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"24", x"6d", x"24", x"00", x"00", x"00", x"00", x"92", x"b6", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"24", x"24", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"00", x"00", x"00", x"b6", x"92", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"00", x"00", x"00", x"b6", x"b6", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"49", x"24", x"24", x"b6", x"b6", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"6d", x"00", x"00", x"00", x"92", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"24", x"00", x"00", x"00", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"6d", x"00", x"00", x"00", x"49", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"b6", x"b6", x"b6", x"92", x"24", x"24", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"00", x"00", x"00", x"00", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"00", x"00", x"00", x"00", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"6d", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"49", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"24", x"6d", x"6d", x"92", x"6d", x"24", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"6d", x"92", x"92", x"92", x"92", x"6d", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"49", x"49", x"49", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"24", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"00", x"00", x"00", x"b6", x"92", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"00", x"00", x"00", x"b6", x"b6", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"49", x"24", x"24", x"b6", x"b6", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"24", x"24", x"24", x"24", x"b6", x"b6", x"b6", x"b6", x"24", x"24", x"24", x"24", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));
	

	constant d_title : memory_m_150_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"00", x"49", x"24", x"db", x"ff", x"ff", x"ff", x"00", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"49", x"b6", x"6d", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"92", x"92", x"b6", x"6d", x"6d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"49", x"49", x"49", x"49", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"ff", x"b6", x"49", x"6d", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"db", x"24", x"92", x"6d", x"6d", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"92", x"49", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"00", x"49", x"24", x"db", x"ff", x"ff", x"ff", x"00", x"49", x"24", x"b6", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"db", x"b6", x"b6", x"b6", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"b6", x"b6", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"b6", x"24", x"49", x"49", x"49", x"49", x"24", x"b6", x"ff", x"ff", x"ff", x"6d", x"49", x"49", x"49", x"92", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"6d", x"6d", x"92", x"92", x"92", x"92", x"6d", x"6d", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"6d", x"49", x"49", x"49", x"49", x"6d", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"db", x"b6", x"b6", x"b6", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"b6", x"b6", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"b6", x"24", x"49", x"49", x"49", x"49", x"24", x"b6", x"ff", x"ff", x"ff", x"6d", x"49", x"49", x"49", x"92", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"6d", x"6d", x"92", x"92", x"92", x"92", x"6d", x"6d", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"6d", x"49", x"49", x"49", x"49", x"6d", x"db", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"49", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"49", x"b6", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"49", x"b6", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"49", x"b6", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"49", x"49", x"49", x"49", x"49", x"49", x"b6", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"49", x"b6", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"49", x"b6", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"49", x"b6", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"6d", x"ff", x"ff", x"ff", x"db", x"24", x"49", x"00", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"db", x"b6", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"b6", x"49", x"92", x"ff", x"ff", x"ff", x"ff", x"b6", x"49", x"6d", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"db", x"24", x"92", x"6d", x"92", x"ff", x"ff", x"db", x"24", x"92", x"6d", x"6d", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"b6", x"49", x"b6", x"92", x"49", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"00", x"49", x"24", x"db", x"ff", x"ff", x"ff", x"00", x"49", x"24", x"b6", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"db", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"b6", x"24", x"49", x"6d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"49", x"92", x"b6", x"00", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"6d", x"6d", x"6d", x"6d", x"49", x"b6", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"b6", x"49", x"b6", x"6d", x"6d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"6d", x"49", x"49", x"49", x"49", x"6d", x"b6", x"92", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"db", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"db", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"92", x"6d", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"92", x"49", x"49", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"ff", x"6d", x"49", x"49", x"49", x"49", x"6d", x"db", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"6d", x"6d", x"92", x"92", x"92", x"92", x"6d", x"6d", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"ff", x"ff", x"ff", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"6d", x"49", x"49", x"49", x"6d", x"ff", x"ff", x"ff", x"b6", x"24", x"49", x"49", x"49", x"49", x"24", x"b6", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"b6", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"db", x"b6", x"b6", x"b6", x"b6", x"db", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"49", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));


	constant d_digit_0 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"6d", x"6d", x"6d", x"6d", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"49", x"6d", x"6d", x"6d", x"6d", x"6d", x"6d", x"49", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));
	
	
	constant d_digit_1 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"24", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));
	
	
	constant d_digit_2 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"24", x"6d", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"49", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"24", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));

	
	constant d_digit_3 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"49", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"6d", x"49", x"24", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"49", x"24", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"49", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"49", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));
	
	
	constant d_digit_4 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"00", x"6d", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"00", x"00", x"00", x"00", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));
	
	
	constant d_digit_5 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"6d", x"49", x"24", x"6d", x"b6", x"b6", x"b6", x"6d", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"92", x"b6", x"6d", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"24", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"49", x"24", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"24", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));
	
	
	constant d_digit_6 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"24", x"49", x"24", x"00", x"00", x"00", x"49", x"49", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"92", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"b6", x"00", x"00", x"00", x"00", x"49", x"6d", x"6d", x"49", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"6d", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"b6", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));

	
	constant d_digit_7 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"24", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));

	
	constant d_digit_8 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"49", x"24", x"24", x"6d", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"6d", x"6d", x"6d", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"92", x"24", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"49", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"00", x"6d", x"b6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"6d", x"6d", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));

	
	constant d_digit_9 : memory_m_20_30 :=
	((x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"6d", x"6d", x"6d", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"b6", x"6d", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"b6", x"b6", x"6d", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"6d", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"b6", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"92", x"24", x"00", x"00", x"00", x"b6", x"24", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"6d", x"b6", x"b6", x"92", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"24", x"00", x"00", x"00", x"92", x"b6", x"b6", x"92", x"24", x"00", x"24", x"b6", x"92", x"6d", x"00", x"00", x"00", x"24", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6d", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"6d", x"49", x"24", x"00", x"00", x"00", x"00", x"24", x"49", x"92", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"), 
	(x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6", x"b6"));
	
	
	constant d_flappy : memory_m_40_40 :=
	((x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"97", x"72", x"6d", x"6d", x"92", x"97", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"04", x"49", x"6d", x"6d", x"24", x"04", x"08", x"76", x"7b", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"29", x"6d", x"ff", x"ff", x"ff", x"fe", x"d9", x"b0", x"24", x"04", x"72", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"97", x"00", x"ff", x"ff", x"ff", x"ff", x"fe", x"fe", x"f9", x"fd", x"d9", x"24", x"28", x"7a", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"5b", x"5b", x"9b", x"6e", x"25", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fe", x"d9", x"fc", x"fd", x"6c", x"00", x"76", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"7b", x"76", x"05", x"00", x"69", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fd", x"d8", x"fc", x"fd", x"90", x"04", x"9b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"76", x"00", x"b2", x"da", x"68", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"d8", x"f8", x"f8", x"fd", x"48", x"24", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"72", x"00", x"da", x"fe", x"d5", x"44", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"f8", x"f5", x"20", x"04", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"00", x"fe", x"fe", x"f9", x"f9", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f8", x"f8", x"f8", x"f9", x"64", x"8c", x"24", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"04", x"b6", x"fe", x"f8", x"f8", x"fd", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f9", x"f8", x"f8", x"f9", x"40", x"f1", x"64", x"4d", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"4d", x"48", x"fe", x"f9", x"d8", x"f8", x"fd", x"44", x"d6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"d9", x"f8", x"f8", x"f9", x"40", x"f0", x"f0", x"20", x"96", x"56", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"00", x"ff", x"fd", x"f8", x"fc", x"fc", x"fc", x"8c", x"8d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f9", x"f8", x"f8", x"f5", x"40", x"f0", x"f0", x"8c", x"49", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"4e", x"48", x"fe", x"f8", x"f8", x"fc", x"f8", x"fc", x"d8", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"d8", x"fc", x"fc", x"ac", x"84", x"f0", x"f0", x"f1", x"20", x"76", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"04", x"da", x"fe", x"f8", x"fc", x"fc", x"f8", x"f8", x"fd", x"44", x"b2", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f8", x"f8", x"f8", x"40", x"f0", x"f0", x"f0", x"f0", x"88", x"4d", x"7b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"97", x"00", x"fe", x"d9", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"d9", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f9", x"f9", x"40", x"cc", x"f0", x"f0", x"f0", x"f0", x"d0", x"24", x"77", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"72", x"28", x"fe", x"d8", x"f8", x"fc", x"f8", x"f8", x"fc", x"f8", x"fc", x"b0", x"20", x"fa", x"ff", x"ff", x"ff", x"ff", x"fd", x"8c", x"20", x"ac", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"20", x"97", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"4d", x"6d", x"fd", x"f8", x"fc", x"f8", x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"d4", x"20", x"68", x"d6", x"fa", x"8d", x"20", x"68", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"44", x"72", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"b1", x"fd", x"f8", x"f8", x"fc", x"fc", x"fc", x"fc", x"f8", x"fc", x"f8", x"fc", x"fd", x"b0", x"68", x"44", x"68", x"f9", x"f9", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"68", x"6d", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"b5", x"fd", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"f8", x"f8", x"fc", x"fc", x"fc", x"fc", x"f8", x"fc", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"88", x"49", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"b5", x"f8", x"f8", x"f8", x"fc", x"fc", x"f8", x"f8", x"fc", x"fd", x"f8", x"f8", x"fd", x"fc", x"f8", x"f8", x"f8", x"fc", x"f8", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"88", x"49", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"28", x"b5", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"fd", x"8c", x"20", x"20", x"24", x"20", x"68", x"d5", x"fc", x"f8", x"fc", x"fc", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"88", x"49", x"7a", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"91", x"fc", x"f8", x"f8", x"f8", x"f8", x"f9", x"20", x"8d", x"ff", x"ff", x"ff", x"ff", x"d6", x"20", x"8c", x"fd", x"fd", x"d4", x"d0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"68", x"4d", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"4d", x"6c", x"fc", x"f8", x"f8", x"fc", x"d9", x"20", x"fa", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"68", x"88", x"60", x"40", x"a4", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"44", x"72", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"72", x"24", x"fd", x"fc", x"f8", x"fd", x"20", x"fb", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"b2", x"40", x"60", x"cd", x"cd", x"80", x"84", x"f0", x"f0", x"f0", x"f0", x"f0", x"24", x"97", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"97", x"00", x"fd", x"f8", x"fd", x"44", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"84", x"ed", x"60", x"cd", x"60", x"cc", x"f0", x"f0", x"f0", x"d0", x"24", x"77", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"28", x"90", x"fd", x"b1", x"44", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"c9", x"e9", x"80", x"cd", x"c9", x"60", x"f0", x"f0", x"f0", x"88", x"4d", x"7b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"52", x"24", x"fe", x"44", x"fb", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"cd", x"ed", x"60", x"cd", x"cd", x"60", x"ec", x"f0", x"f1", x"20", x"76", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7a", x"04", x"d6", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"f1", x"e8", x"60", x"cd", x"c9", x"a4", x"a8", x"f1", x"8c", x"49", x"76", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"72", x"00", x"44", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"40", x"f6", x"ed", x"60", x"cd", x"c9", x"a4", x"84", x"d1", x"24", x"97", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"40", x"f6", x"ed", x"60", x"cd", x"e9", x"c8", x"84", x"24", x"76", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"04", x"92", x"ff", x"ff", x"ff", x"ff", x"fb", x"b2", x"d6", x"ff", x"ff", x"ff", x"ff", x"20", x"f6", x"f1", x"60", x"c9", x"e9", x"c9", x"20", x"72", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"96", x"00", x"b7", x"ff", x"ff", x"92", x"20", x"20", x"20", x"20", x"d7", x"ff", x"ff", x"40", x"f6", x"f1", x"60", x"cd", x"e9", x"a8", x"49", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"77", x"00", x"6e", x"ff", x"8e", x"20", x"44", x"45", x"20", x"20", x"ff", x"ff", x"40", x"f6", x"f1", x"60", x"e9", x"e9", x"a8", x"49", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"9b", x"29", x"00", x"d7", x"92", x"ff", x"ff", x"8e", x"d7", x"ff", x"d6", x"40", x"f6", x"f1", x"80", x"c9", x"e9", x"88", x"4d", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"76", x"09", x"00", x"49", x"92", x"b6", x"b2", x"69", x"20", x"20", x"f6", x"ed", x"80", x"ed", x"e9", x"84", x"4d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"97", x"72", x"4d", x"29", x"29", x"49", x"6d", x"20", x"f1", x"ed", x"80", x"cd", x"ed", x"40", x"76", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"5b", x"7b", x"77", x"7b", x"97", x"25", x"d1", x"ed", x"60", x"cd", x"cd", x"20", x"97", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"29", x"ad", x"c9", x"40", x"69", x"65", x"49", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"72", x"20", x"44", x"6e", x"29", x"29", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"6d", x"6d", x"97", x"77", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"));
	
	
	constant d_flappy_bg_status : memory_m_40_40_bg :=
	(('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'));
	
	
	constant d_flappy_incr : memory_m_40_40 :=
	((x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"77", x"7b", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"4e", x"04", x"04", x"4d", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"77", x"7b", x"7b", x"77", x"76", x"77", x"7b", x"05", x"25", x"fb", x"fb", x"49", x"04", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"72", x"29", x"04", x"00", x"24", x"24", x"24", x"00", x"8e", x"ff", x"ff", x"ff", x"ff", x"6d", x"04", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"52", x"04", x"04", x"91", x"fa", x"ff", x"ff", x"ff", x"b1", x"44", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"48", x"29", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"77", x"24", x"24", x"da", x"fe", x"fe", x"fd", x"fd", x"f9", x"fa", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fe", x"04", x"76", x"77", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"76", x"00", x"91", x"fe", x"fe", x"f9", x"d8", x"d8", x"f8", x"fc", x"68", x"8d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"d9", x"d9", x"04", x"7a", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"52", x"00", x"fa", x"fe", x"f9", x"f8", x"f8", x"fc", x"f8", x"f8", x"f9", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f9", x"fd", x"6c", x"51", x"77", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"76", x"00", x"fe", x"fe", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"90", x"68", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fd", x"f8", x"f9", x"04", x"7b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"00", x"fe", x"fd", x"f8", x"f8", x"f8", x"f8", x"fc", x"fc", x"f8", x"fd", x"20", x"fa", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f9", x"f8", x"fd", x"28", x"72", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"04", x"b5", x"fd", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"f9", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"d9", x"d8", x"fc", x"8c", x"4d", x"7b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"4d", x"48", x"fd", x"f8", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"b0", x"48", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"d8", x"fc", x"f8", x"b1", x"49", x"7a", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"00", x"fe", x"f8", x"fc", x"fc", x"f8", x"f8", x"f8", x"f8", x"fc", x"f8", x"f8", x"b0", x"68", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"fc", x"b1", x"48", x"7a", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"2d", x"6c", x"fd", x"f8", x"f8", x"fc", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"fc", x"b0", x"44", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f8", x"f8", x"f8", x"fc", x"8c", x"00", x"7b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"97", x"04", x"d9", x"f8", x"fc", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"f8", x"fc", x"f8", x"f9", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f9", x"f8", x"f8", x"f8", x"f9", x"44", x"44", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"72", x"24", x"fd", x"fc", x"fc", x"f8", x"f8", x"fc", x"f8", x"fc", x"fc", x"f8", x"f8", x"f8", x"fd", x"48", x"b1", x"ff", x"ff", x"ff", x"ff", x"fe", x"fd", x"d8", x"f8", x"f8", x"fd", x"44", x"cc", x"64", x"72", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7a", x"4d", x"8c", x"fd", x"fc", x"fc", x"fd", x"d4", x"8c", x"8c", x"8c", x"b0", x"f8", x"fc", x"f8", x"f8", x"d8", x"20", x"ff", x"ff", x"ff", x"fe", x"f9", x"d8", x"fc", x"f8", x"fd", x"88", x"64", x"f1", x"68", x"72", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7a", x"24", x"d5", x"fd", x"d5", x"48", x"20", x"48", x"91", x"b6", x"b6", x"8d", x"20", x"68", x"fd", x"f8", x"fc", x"b0", x"20", x"d6", x"fa", x"fa", x"fe", x"fd", x"fd", x"d5", x"64", x"60", x"f0", x"f0", x"88", x"52", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7a", x"04", x"fa", x"68", x"20", x"d6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"8d", x"44", x"fd", x"f8", x"fc", x"d4", x"44", x"20", x"20", x"40", x"44", x"40", x"40", x"a8", x"f0", x"f0", x"f0", x"64", x"72", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"24", x"64", x"8d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"6c", x"6c", x"fc", x"f8", x"fc", x"fc", x"fd", x"f9", x"d0", x"d0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"44", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"00", x"69", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"f9", x"f8", x"fc", x"fc", x"f8", x"f4", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"40", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"00", x"f7", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"68", x"8c", x"fc", x"f8", x"f8", x"f8", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"d1", x"44", x"7a", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"00", x"fb", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"89", x"64", x"fd", x"fc", x"f8", x"d0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"68", x"6d", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"05", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"40", x"40", x"60", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"20", x"97", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"4d", x"92", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"d6", x"20", x"60", x"cd", x"a8", x"60", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ac", x"29", x"77", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"76", x"25", x"ff", x"fb", x"8d", x"d6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"40", x"80", x"e9", x"c9", x"c9", x"60", x"f1", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f1", x"20", x"76", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"05", x"ff", x"24", x"20", x"20", x"69", x"ff", x"ff", x"ff", x"ff", x"ff", x"69", x"64", x"ed", x"e9", x"80", x"c8", x"80", x"cc", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"68", x"49", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"52", x"25", x"8e", x"45", x"20", x"20", x"8e", x"ff", x"ff", x"ff", x"d6", x"40", x"f2", x"c9", x"a4", x"a0", x"ed", x"80", x"cc", x"f0", x"f0", x"f0", x"f0", x"f0", x"ac", x"00", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"92", x"ff", x"fb", x"20", x"20", x"ff", x"ff", x"ff", x"20", x"f6", x"f1", x"c9", x"60", x"ed", x"ec", x"60", x"cc", x"f0", x"f0", x"f0", x"f0", x"d1", x"20", x"76", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"77", x"04", x"b6", x"ff", x"20", x"69", x"ff", x"ff", x"40", x"cd", x"f2", x"cd", x"60", x"c9", x"e9", x"e8", x"60", x"f1", x"f0", x"f0", x"f0", x"d0", x"00", x"76", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"00", x"6d", x"ff", x"ff", x"ff", x"8d", x"64", x"f6", x"f1", x"84", x"a4", x"ed", x"e9", x"a4", x"a8", x"f0", x"f0", x"f1", x"8c", x"20", x"76", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"77", x"29", x"00", x"6d", x"69", x"40", x"f6", x"f1", x"a8", x"60", x"ed", x"c9", x"cd", x"60", x"f0", x"f0", x"d1", x"44", x"29", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"72", x"24", x"20", x"cd", x"f2", x"ed", x"60", x"e9", x"e8", x"cd", x"64", x"88", x"ac", x"64", x"44", x"72", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"96", x"40", x"f6", x"f1", x"80", x"c4", x"e9", x"e9", x"a9", x"20", x"29", x"4d", x"76", x"7a", x"76", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"25", x"d1", x"ed", x"a8", x"80", x"e9", x"e9", x"cd", x"20", x"96", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"96", x"20", x"f2", x"c9", x"80", x"ed", x"e8", x"cd", x"20", x"72", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"4e", x"49", x"89", x"40", x"a4", x"cd", x"cd", x"40", x"72", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"09", x"29", x"49", x"89", x"89", x"20", x"72", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"77", x"96", x"44", x"64", x"92", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"));
	
	
	constant d_flappy_incr_bg_status : memory_m_40_40_bg :=
	(('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'));

	
	constant d_flappy_decr : memory_m_40_40 :=
	((x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"76", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"77", x"97", x"96", x"72", x"72", x"72", x"77", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"7b", x"56", x"2d", x"04", x"00", x"24", x"48", x"48", x"28", x"00", x"28", x"51", x"56", x"76", x"7b", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"72", x"00", x"24", x"91", x"d9", x"fd", x"fd", x"fc", x"fc", x"fc", x"fd", x"b4", x"44", x"20", x"24", x"24", x"6d", x"77", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"52", x"00", x"fb", x"fe", x"fe", x"fe", x"fd", x"fc", x"f8", x"f8", x"f8", x"fc", x"f8", x"fd", x"88", x"ac", x"d1", x"68", x"24", x"4d", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"04", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fe", x"fd", x"d8", x"f8", x"f8", x"f8", x"fd", x"40", x"d1", x"f0", x"d0", x"88", x"20", x"76", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"76", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fd", x"f8", x"f8", x"f8", x"f8", x"d0", x"40", x"f0", x"f0", x"f0", x"d1", x"00", x"72", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"f8", x"fd", x"40", x"cc", x"f0", x"f0", x"f0", x"f1", x"20", x"71", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"29", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fd", x"f8", x"f8", x"f9", x"88", x"a8", x"f0", x"f0", x"f0", x"ec", x"f1", x"20", x"72", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"97", x"29", x"00", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f8", x"f8", x"f9", x"8c", x"a8", x"f0", x"f0", x"f0", x"f0", x"f0", x"d1", x"20", x"76", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"72", x"24", x"6d", x"6d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f9", x"68", x"cc", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"d0", x"00", x"97", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"b6", x"fe", x"20", x"b6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f9", x"f9", x"40", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"68", x"4d", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"00", x"ff", x"f9", x"f9", x"20", x"d6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f9", x"8c", x"64", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"d1", x"20", x"76", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"52", x"49", x"ff", x"f8", x"f8", x"d8", x"20", x"da", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fa", x"20", x"f9", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"88", x"4d", x"7b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"77", x"2d", x"6d", x"fe", x"f8", x"f8", x"fc", x"d9", x"20", x"b1", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"24", x"90", x"fd", x"f4", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"d0", x"24", x"77", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"77", x"29", x"96", x"fe", x"f8", x"f8", x"f8", x"f8", x"f9", x"24", x"24", x"d6", x"ff", x"ff", x"ff", x"da", x"44", x"44", x"fd", x"f8", x"f8", x"d0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"24", x"96", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"7b", x"09", x"b6", x"fe", x"f8", x"fc", x"f8", x"f8", x"f8", x"fd", x"b0", x"44", x"20", x"20", x"20", x"20", x"b0", x"fd", x"f8", x"f8", x"f8", x"f4", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"68", x"72", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"7b", x"29", x"b5", x"fe", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"fc", x"f8", x"fd", x"fc", x"fc", x"f8", x"f8", x"fc", x"f8", x"f9", x"88", x"84", x"a8", x"ec", x"f0", x"f0", x"f0", x"f0", x"8c", x"6d", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"77", x"2d", x"91", x"fe", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"fc", x"fc", x"f8", x"fc", x"f8", x"fc", x"fc", x"fc", x"fd", x"fd", x"64", x"84", x"a8", x"84", x"60", x"60", x"f0", x"f0", x"f0", x"ad", x"49", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"52", x"49", x"fe", x"f8", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"fc", x"fc", x"fd", x"d4", x"68", x"44", x"44", x"44", x"8d", x"40", x"cd", x"c4", x"a4", x"cd", x"a8", x"60", x"cc", x"f1", x"b1", x"48", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"00", x"fe", x"f8", x"f8", x"fc", x"f8", x"fc", x"f8", x"fc", x"f8", x"f8", x"fd", x"44", x"44", x"d6", x"fb", x"fb", x"8d", x"20", x"40", x"c8", x"ed", x"60", x"c9", x"cd", x"c9", x"60", x"d1", x"ad", x"6d", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"00", x"fe", x"f9", x"fc", x"f8", x"f8", x"f8", x"fc", x"f8", x"f8", x"fd", x"20", x"d6", x"ff", x"ff", x"ff", x"ff", x"ff", x"fb", x"20", x"84", x"c9", x"c9", x"80", x"e9", x"e9", x"c8", x"40", x"8d", x"6d", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"49", x"8d", x"fd", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"68", x"b1", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"d6", x"40", x"cd", x"cd", x"80", x"c4", x"e9", x"e9", x"a4", x"20", x"92", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"96", x"00", x"fe", x"d8", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"64", x"ad", x"f1", x"cd", x"60", x"ed", x"e9", x"ed", x"40", x"92", x"76", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"28", x"91", x"fd", x"fc", x"fc", x"f8", x"f8", x"fc", x"90", x"8d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"f6", x"f1", x"a4", x"80", x"e9", x"e9", x"a9", x"44", x"7b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"00", x"fe", x"f8", x"f8", x"fc", x"f8", x"f9", x"68", x"da", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"89", x"88", x"f1", x"ed", x"60", x"c8", x"e9", x"ed", x"40", x"72", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"4d", x"48", x"fd", x"f8", x"f8", x"f8", x"fd", x"40", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"20", x"f2", x"f5", x"cd", x"60", x"e9", x"e8", x"a9", x"25", x"77", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"04", x"90", x"f9", x"f8", x"f8", x"fd", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"d6", x"40", x"f6", x"f1", x"84", x"a4", x"e8", x"cd", x"20", x"97", x"77", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"00", x"b5", x"fd", x"f8", x"fd", x"20", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"44", x"ad", x"f6", x"cd", x"60", x"ed", x"c9", x"65", x"6e", x"77", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"7b", x"76", x"04", x"90", x"fd", x"fd", x"24", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fb", x"44", x"20", x"20", x"b2", x"ff", x"b2", x"20", x"f2", x"f1", x"c8", x"80", x"cd", x"69", x"4d", x"77", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"76", x"04", x"68", x"fe", x"68", x"d6", x"ff", x"ff", x"ff", x"ff", x"ff", x"db", x"20", x"20", x"20", x"20", x"89", x"ff", x"24", x"20", x"40", x"f6", x"cd", x"60", x"40", x"20", x"72", x"77", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5a", x"7a", x"2d", x"00", x"8d", x"40", x"ff", x"ff", x"ff", x"ff", x"ff", x"69", x"20", x"44", x"ff", x"ff", x"ff", x"24", x"04", x"96", x"4d", x"44", x"d2", x"64", x"8e", x"72", x"77", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"77", x"96", x"25", x"00", x"24", x"db", x"ff", x"ff", x"ff", x"ff", x"69", x"b6", x"ff", x"6e", x"00", x"4d", x"97", x"5b", x"77", x"4d", x"24", x"04", x"72", x"77", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"56", x"7b", x"76", x"2d", x"04", x"04", x"49", x"4d", x"6d", x"49", x"04", x"04", x"2e", x"77", x"77", x"5b", x"5b", x"5b", x"7b", x"52", x"32", x"7b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5a", x"5a", x"5b", x"77", x"7b", x"76", x"72", x"72", x"72", x"72", x"77", x"7b", x"7b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"77", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"));

	
	constant d_flappy_decr_bg_status : memory_m_40_40_bg :=
	(('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '1', '1', '1', '1', '1', '1', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '1', '1', '1', '1', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'), 
	('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'));
	
	
	constant d_flappy_dead : memory_m_40_40 :=
	((x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"29", x"2a", x"32", x"5b", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"65", x"8d", x"88", x"64", x"45", x"25", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"64", x"ff", x"ff", x"ff", x"fc", x"d4", x"ac", x"60", x"21", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"d6", x"ff", x"ff", x"ff", x"ff", x"fe", x"fc", x"fc", x"d0", x"64", x"25", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"2e", x"65", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fc", x"fc", x"fc", x"88", x"21", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"25", x"20", x"89", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"fc", x"fc", x"a8", x"21", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"36", x"20", x"ad", x"b2", x"69", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"f8", x"f8", x"fc", x"fc", x"84", x"21", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"36", x"20", x"d2", x"ff", x"d4", x"65", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"fc", x"d8", x"40", x"21", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"d2", x"ff", x"fc", x"d4", x"40", x"fb", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"f8", x"f8", x"fc", x"f8", x"a8", x"a0", x"25", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"a9", x"ff", x"fc", x"fc", x"f8", x"40", x"b7", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"f8", x"fc", x"f8", x"88", x"f0", x"80", x"2a", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"2e", x"60", x"ff", x"fd", x"f8", x"fc", x"fc", x"64", x"8e", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"fc", x"d8", x"64", x"ec", x"f0", x"40", x"37", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"d6", x"fe", x"f8", x"f8", x"f8", x"fc", x"88", x"65", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"f8", x"fc", x"d4", x"60", x"ec", x"f4", x"c8", x"29", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"64", x"ff", x"fc", x"f8", x"f8", x"f8", x"fc", x"d4", x"41", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"f8", x"fc", x"8c", x"40", x"f0", x"f0", x"f0", x"64", x"37", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"ad", x"fe", x"f8", x"f8", x"f8", x"fc", x"fc", x"fc", x"44", x"8e", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f8", x"fc", x"f8", x"20", x"c8", x"f0", x"f0", x"f0", x"a4", x"2a", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"40", x"da", x"fd", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"d4", x"20", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"fc", x"fc", x"20", x"84", x"f4", x"f0", x"f0", x"f0", x"ec", x"45", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"65", x"fe", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"8c", x"20", x"b7", x"ff", x"ff", x"ff", x"ff", x"fc", x"8c", x"20", x"84", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"64", x"37", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2a", x"89", x"fe", x"f8", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"fc", x"b0", x"20", x"66", x"b3", x"d7", x"8e", x"40", x"40", x"ac", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"84", x"2e", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"ad", x"fd", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"fc", x"f8", x"88", x"44", x"40", x"64", x"b0", x"fc", x"f4", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"a4", x"2a", x"5f", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"ad", x"fd", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"f8", x"fc", x"fc", x"fc", x"f0", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"c8", x"29", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"ad", x"fc", x"f8", x"f8", x"fc", x"fc", x"f8", x"fc", x"fc", x"fc", x"d4", x"b4", x"d8", x"fc", x"fc", x"fc", x"fc", x"f8", x"fc", x"f4", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"c8", x"29", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"ac", x"fc", x"f8", x"f8", x"fc", x"f8", x"fc", x"fc", x"8c", x"44", x"65", x"65", x"64", x"64", x"d4", x"fc", x"fc", x"fc", x"fc", x"f4", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"c8", x"29", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"ac", x"fc", x"fc", x"f8", x"f8", x"fc", x"f8", x"40", x"65", x"d7", x"ff", x"ff", x"fb", x"8e", x"41", x"68", x"fc", x"fc", x"b4", x"cc", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"a4", x"29", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"88", x"fc", x"fc", x"f8", x"fc", x"f8", x"20", x"b3", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"21", x"68", x"8c", x"40", x"40", x"84", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"84", x"2e", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"64", x"fc", x"fc", x"fc", x"fc", x"40", x"d7", x"df", x"b6", x"ff", x"ff", x"ff", x"ff", x"b6", x"ff", x"d6", x"00", x"20", x"e8", x"e8", x"40", x"64", x"f0", x"f0", x"f0", x"f0", x"f0", x"64", x"32", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"40", x"d4", x"fc", x"fc", x"64", x"8e", x"db", x"00", x"00", x"d7", x"ff", x"ff", x"6d", x"00", x"49", x"ff", x"41", x"80", x"ec", x"a4", x"e8", x"40", x"88", x"f0", x"f0", x"f0", x"ec", x"45", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"25", x"8c", x"fc", x"b0", x"69", x"b6", x"00", x"00", x"00", x"00", x"ff", x"92", x"00", x"00", x"00", x"24", x"45", x"a4", x"ec", x"60", x"e8", x"c8", x"40", x"f0", x"f0", x"f0", x"a4", x"29", x"5f", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"64", x"fc", x"64", x"b3", x"ff", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"65", x"c4", x"e8", x"84", x"c8", x"ec", x"60", x"ac", x"f0", x"f0", x"64", x"33", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"45", x"88", x"88", x"ff", x"ff", x"d6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"ff", x"89", x"ed", x"e8", x"84", x"c8", x"ec", x"84", x"88", x"f4", x"c8", x"29", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"52", x"20", x"65", x"ff", x"ff", x"ff", x"b6", x"00", x"00", x"00", x"00", x"00", x"49", x"ff", x"ff", x"69", x"f1", x"ec", x"80", x"c8", x"ec", x"a4", x"88", x"f0", x"60", x"37", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"40", x"ff", x"ff", x"ff", x"6d", x"00", x"00", x"00", x"00", x"00", x"24", x"ff", x"ff", x"65", x"f1", x"ed", x"80", x"c8", x"ec", x"a4", x"84", x"84", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"ad", x"ff", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"db", x"89", x"f1", x"f1", x"80", x"c8", x"ec", x"c8", x"20", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"65", x"40", x"00", x"00", x"00", x"00", x"49", x"00", x"00", x"00", x"00", x"00", x"89", x"f1", x"f1", x"80", x"c8", x"ec", x"c4", x"25", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"20", x"00", x"00", x"00", x"6d", x"ff", x"b6", x"00", x"00", x"00", x"4d", x"89", x"f1", x"f1", x"80", x"c8", x"ec", x"c4", x"29", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"49", x"00", x"20", x"ff", x"ff", x"ff", x"b6", x"00", x"b6", x"fb", x"40", x"f1", x"f1", x"84", x"c8", x"ec", x"c0", x"29", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"49", x"65", x"89", x"b2", x"f7", x"ae", x"ae", x"40", x"40", x"f1", x"f1", x"a4", x"c8", x"ec", x"a0", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"36", x"2d", x"25", x"25", x"45", x"25", x"29", x"45", x"ed", x"f1", x"a4", x"c8", x"ec", x"80", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"c8", x"ed", x"84", x"c8", x"e8", x"64", x"37", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"c4", x"ed", x"20", x"a0", x"c0", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"80", x"80", x"29", x"49", x"45", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"));
	
	
	constant d_flappy_dead_incr : memory_m_40_40 :=
	((x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"2e", x"20", x"20", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"5b", x"32", x"32", x"5b", x"5b", x"25", x"60", x"d6", x"d6", x"64", x"21", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"29", x"25", x"45", x"45", x"65", x"69", x"20", x"65", x"ff", x"ff", x"ff", x"ff", x"84", x"21", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"32", x"20", x"40", x"8d", x"d6", x"fb", x"ff", x"ff", x"8d", x"40", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"84", x"25", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"25", x"40", x"ad", x"ff", x"ff", x"fe", x"fd", x"fc", x"fc", x"40", x"b7", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fc", x"40", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"20", x"89", x"ff", x"ff", x"fd", x"f8", x"f8", x"f8", x"fc", x"68", x"65", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"d4", x"25", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"32", x"20", x"b2", x"ff", x"fd", x"f8", x"f8", x"f8", x"fc", x"fc", x"f8", x"40", x"d7", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"fc", x"88", x"2a", x"5f", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"36", x"20", x"d2", x"fe", x"fc", x"f8", x"f8", x"fc", x"f8", x"f8", x"fc", x"8c", x"45", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"fc", x"f8", x"45", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"b2", x"fe", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"fc", x"44", x"92", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"fc", x"88", x"2e", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"25", x"89", x"fd", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"d4", x"40", x"db", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"f8", x"fc", x"ac", x"29", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"2e", x"60", x"fd", x"fc", x"f8", x"f8", x"f8", x"fc", x"f8", x"f8", x"f8", x"fc", x"b0", x"65", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"f8", x"fc", x"fc", x"d0", x"29", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"21", x"d5", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"8c", x"69", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f8", x"f8", x"fc", x"d0", x"25", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"2e", x"84", x"fc", x"f8", x"fc", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"b0", x"65", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"f8", x"f8", x"fc", x"ac", x"21", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"d0", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"d8", x"40", x"fb", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"fc", x"fc", x"64", x"60", x"32", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"44", x"fc", x"fc", x"f8", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"f8", x"f8", x"fc", x"64", x"8e", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"fc", x"fc", x"68", x"a4", x"a8", x"2e", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"2a", x"88", x"fc", x"fc", x"fc", x"fc", x"b0", x"8c", x"68", x"68", x"8c", x"d8", x"fc", x"fc", x"fc", x"d4", x"20", x"db", x"ff", x"ff", x"ff", x"fd", x"f8", x"fc", x"fc", x"fc", x"6c", x"40", x"f4", x"a8", x"2e", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"b0", x"fc", x"d4", x"88", x"8d", x"ae", x"b2", x"8e", x"8e", x"8a", x"45", x"68", x"fc", x"fc", x"fc", x"b0", x"21", x"8f", x"da", x"f8", x"fc", x"fc", x"fc", x"d4", x"44", x"40", x"ec", x"f4", x"a4", x"2e", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"45", x"f4", x"8c", x"41", x"6a", x"8e", x"72", x"b6", x"ff", x"ff", x"ff", x"ff", x"66", x"44", x"fc", x"fc", x"fc", x"b0", x"40", x"64", x"64", x"44", x"64", x"64", x"40", x"80", x"f0", x"f0", x"f0", x"a4", x"2e", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"69", x"60", x"65", x"ff", x"71", x"00", x"00", x"00", x"db", x"ff", x"ff", x"ff", x"ff", x"6a", x"68", x"fc", x"f8", x"fc", x"fc", x"fc", x"d4", x"a8", x"a4", x"cc", x"f0", x"f0", x"f0", x"f0", x"f0", x"84", x"32", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"41", x"ff", x"ff", x"6d", x"00", x"00", x"00", x"92", x"ff", x"ff", x"ff", x"ff", x"ff", x"40", x"d4", x"fc", x"f8", x"fc", x"fc", x"f8", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"64", x"37", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"b2", x"ff", x"ff", x"b6", x"00", x"00", x"00", x"6d", x"ff", x"db", x"92", x"b6", x"ff", x"6a", x"68", x"fc", x"fc", x"fc", x"f8", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ec", x"49", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"d2", x"ff", x"ff", x"db", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"24", x"ff", x"8e", x"44", x"fc", x"fc", x"fc", x"f0", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"a8", x"2e", x"5f", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"49", x"89", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"df", x"89", x"20", x"64", x"68", x"d0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"64", x"33", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"52", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"20", x"40", x"e4", x"80", x"40", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4", x"c8", x"25", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6d", x"bb", x"49", x"40", x"ec", x"ec", x"c8", x"60", x"cc", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"60", x"32", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"6d", x"ff", x"ff", x"92", x"40", x"ec", x"ec", x"60", x"a4", x"84", x"a8", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4", x"a4", x"25", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"20", x"db", x"ff", x"db", x"00", x"00", x"00", x"49", x"ff", x"b6", x"40", x"f1", x"ec", x"84", x"60", x"ec", x"80", x"a8", x"f0", x"f0", x"f0", x"f0", x"f4", x"c8", x"20", x"37", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"49", x"ae", x"ff", x"ff", x"00", x"00", x"00", x"24", x"db", x"40", x"cd", x"f5", x"c4", x"40", x"e8", x"ec", x"60", x"ac", x"f0", x"f0", x"f0", x"f4", x"ec", x"40", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"ae", x"ff", x"49", x"00", x"00", x"24", x"45", x"a8", x"f9", x"ec", x"40", x"a4", x"ec", x"e8", x"40", x"ec", x"f0", x"f0", x"f4", x"ec", x"40", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"a9", x"db", x"96", x"df", x"6d", x"60", x"f5", x"f1", x"80", x"60", x"ec", x"ec", x"84", x"64", x"f0", x"f0", x"f4", x"c8", x"40", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"60", x"d6", x"b2", x"40", x"d1", x"f9", x"c8", x"40", x"e8", x"e8", x"e8", x"60", x"cc", x"f4", x"ec", x"a4", x"25", x"37", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"4e", x"20", x"00", x"a9", x"fa", x"ed", x"40", x"a4", x"ec", x"ec", x"80", x"64", x"ec", x"84", x"45", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"37", x"40", x"f5", x"f1", x"80", x"84", x"ec", x"ec", x"c4", x"20", x"45", x"49", x"32", x"3b", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"a8", x"f5", x"c4", x"60", x"e8", x"ec", x"e8", x"40", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"37", x"65", x"f1", x"e8", x"60", x"c8", x"ec", x"e8", x"60", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"a0", x"e4", x"20", x"84", x"ec", x"e8", x"80", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"45", x"29", x"05", x"c0", x"e4", x"60", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"45", x"45", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"));
	
	
	constant d_flappy_dead_decr : memory_m_40_40 :=
	((x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"5b", x"37", x"33", x"32", x"33", x"5b", x"5b", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"2a", x"25", x"45", x"68", x"68", x"68", x"68", x"45", x"25", x"2e", x"5b", x"37", x"5b", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"36", x"20", x"60", x"88", x"d0", x"f4", x"f8", x"fc", x"fc", x"fc", x"f8", x"ac", x"60", x"20", x"64", x"49", x"2e", x"3b", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"20", x"d1", x"fe", x"fe", x"fe", x"fd", x"fc", x"f8", x"f8", x"fc", x"fc", x"fc", x"fc", x"68", x"80", x"ec", x"84", x"40", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"d2", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fc", x"f8", x"f8", x"f8", x"fc", x"fc", x"40", x"cc", x"f4", x"ec", x"80", x"25", x"37", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"45", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"f8", x"fc", x"b0", x"40", x"f0", x"f0", x"f4", x"e8", x"40", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"45", x"d6", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"f8", x"f8", x"fc", x"fc", x"44", x"a8", x"f0", x"f0", x"f4", x"ec", x"60", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"8d", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"f8", x"fc", x"68", x"84", x"f0", x"f0", x"f0", x"f0", x"f0", x"60", x"2e", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"40", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"f8", x"fc", x"68", x"84", x"f0", x"f0", x"f0", x"f0", x"f0", x"ec", x"40", x"33", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"69", x"65", x"69", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fd", x"f8", x"fc", x"68", x"84", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4", x"c8", x"20", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"b1", x"fe", x"20", x"8e", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fe", x"fc", x"fc", x"44", x"c8", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4", x"84", x"2a", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"45", x"fb", x"fd", x"d8", x"20", x"b2", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"fc", x"90", x"40", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"40", x"37", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"65", x"ff", x"fc", x"fc", x"d4", x"20", x"b2", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"f9", x"20", x"b0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f4", x"84", x"2a", x"5f", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"89", x"ff", x"fc", x"f8", x"fc", x"d4", x"00", x"8e", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"45", x"68", x"fc", x"f4", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"ec", x"45", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"89", x"fe", x"f8", x"f8", x"f8", x"fc", x"d8", x"40", x"41", x"b6", x"fb", x"ff", x"ff", x"db", x"45", x"40", x"fc", x"fc", x"fc", x"f0", x"ec", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"64", x"32", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"ad", x"fe", x"f8", x"f8", x"f8", x"f8", x"fc", x"fc", x"8c", x"40", x"40", x"41", x"40", x"40", x"68", x"fc", x"fc", x"f8", x"fc", x"f8", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"f0", x"a4", x"2e", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5f", x"25", x"ad", x"fe", x"f8", x"fc", x"fc", x"f8", x"f8", x"fc", x"fc", x"fc", x"d4", x"b4", x"d4", x"f8", x"fc", x"fc", x"f8", x"fc", x"fc", x"fc", x"88", x"64", x"88", x"cc", x"f0", x"f0", x"f0", x"f0", x"c8", x"2e", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"89", x"fe", x"f8", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"fc", x"8c", x"40", x"84", x"80", x"60", x"64", x"cc", x"f0", x"f0", x"e8", x"49", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"65", x"fe", x"fc", x"f8", x"f8", x"f8", x"f8", x"fc", x"fc", x"f8", x"f8", x"fc", x"fc", x"b4", x"68", x"64", x"64", x"64", x"8c", x"40", x"e8", x"e8", x"a4", x"ec", x"80", x"20", x"ac", x"f4", x"e8", x"49", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"65", x"fe", x"fc", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"f8", x"fc", x"fc", x"64", x"45", x"8e", x"b3", x"d7", x"8e", x"00", x"20", x"c8", x"e8", x"40", x"c8", x"ec", x"c4", x"20", x"cc", x"ec", x"49", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"24", x"d6", x"fd", x"f8", x"f8", x"f8", x"fc", x"f8", x"f8", x"fc", x"fc", x"40", x"66", x"ff", x"ff", x"ff", x"df", x"ff", x"fb", x"20", x"60", x"ec", x"a4", x"40", x"e8", x"ec", x"c4", x"40", x"c8", x"4e", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"89", x"fe", x"f8", x"f8", x"f8", x"f8", x"f8", x"f8", x"fc", x"88", x"66", x"ff", x"ff", x"ff", x"db", x"00", x"00", x"49", x"6d", x"40", x"e8", x"ec", x"60", x"84", x"ec", x"ec", x"a4", x"20", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"40", x"fa", x"fc", x"f8", x"f8", x"fc", x"f8", x"fc", x"d8", x"65", x"ff", x"ff", x"ff", x"ff", x"92", x"00", x"00", x"00", x"92", x"8e", x"88", x"f5", x"c4", x"40", x"c8", x"e8", x"e8", x"60", x"32", x"5f", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"25", x"8d", x"fd", x"f8", x"f8", x"f8", x"f8", x"fc", x"8c", x"69", x"b6", x"92", x"ff", x"ff", x"49", x"00", x"00", x"00", x"df", x"ff", x"40", x"f1", x"f1", x"80", x"60", x"ec", x"ec", x"c4", x"25", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"41", x"f9", x"fc", x"f8", x"f8", x"fc", x"fc", x"ac", x"45", x"00", x"00", x"00", x"49", x"00", x"00", x"00", x"24", x"ff", x"ff", x"69", x"64", x"fa", x"ed", x"60", x"a4", x"ec", x"e8", x"80", x"32", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"29", x"64", x"fd", x"fc", x"f8", x"fc", x"fc", x"88", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"db", x"ff", x"ff", x"45", x"cd", x"f9", x"c8", x"40", x"e8", x"ec", x"c4", x"25", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"21", x"ac", x"fc", x"fc", x"fc", x"fc", x"68", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"8e", x"60", x"f5", x"f1", x"80", x"84", x"ec", x"e8", x"64", x"36", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"20", x"ac", x"fc", x"fc", x"f8", x"64", x"db", x"b6", x"49", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"b6", x"8e", x"88", x"f9", x"ed", x"60", x"c8", x"ec", x"a0", x"2e", x"5f", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"20", x"ac", x"fc", x"fc", x"44", x"d7", x"ff", x"ff", x"b6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ff", x"b6", x"00", x"d1", x"f5", x"a4", x"60", x"ec", x"c4", x"29", x"5f", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"21", x"84", x"fc", x"8c", x"8e", x"ff", x"ff", x"91", x"00", x"00", x"00", x"6d", x"b6", x"49", x"00", x"6d", x"ff", x"69", x"00", x"64", x"f1", x"ed", x"60", x"60", x"80", x"52", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"60", x"88", x"44", x"ff", x"ff", x"24", x"00", x"00", x"00", x"db", x"ff", x"ff", x"ff", x"ff", x"85", x"20", x"5b", x"2e", x"60", x"f1", x"a4", x"09", x"36", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"32", x"45", x"20", x"64", x"d6", x"00", x"00", x"00", x"24", x"ff", x"ff", x"fb", x"d2", x"40", x"25", x"5b", x"5f", x"5b", x"2e", x"80", x"80", x"36", x"5f", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"25", x"20", x"40", x"20", x"00", x"45", x"ae", x"69", x"45", x"25", x"32", x"5f", x"5b", x"5b", x"5b", x"5b", x"2e", x"29", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"5b", x"52", x"52", x"4e", x"2d", x"32", x"5b", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5f", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"));
	
	
	constant d_start_game_text : memory_m_255_30 :=
	((x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"32", x"2d", x"09", x"09", x"09", x"09", x"2d", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"09", x"09", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"52", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"04", x"00", x"00", x"00", x"05", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"04", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"2e", x"29", x"00", x"00", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"56", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"32", x"32", x"5b", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"2d", x"2d", x"5b", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"09", x"00", x"00", x"00", x"00", x"09", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"05", x"32", x"5b", x"5b", x"5b", x"5b", x"56", x"08", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"04", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"05", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"29", x"00", x"00", x"00", x"00", x"00", x"04", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2e", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"2d", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"56", x"2d", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"2d", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"09", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"29", x"00", x"00", x"00", x"00", x"09", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"09", x"5b", x"00", x"00", x"00", x"5b", x"32", x"04", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"56", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"09", x"56", x"00", x"00", x"00", x"5b", x"5b", x"09", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"2d", x"09", x"04", x"04", x"5b", x"5b", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"32", x"32", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"2e", x"00", x"00", x"00", x"00", x"2e", x"2e", x"2e", x"32", x"2e", x"32", x"2e", x"32", x"2e", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"2d", x"00", x"00", x"00", x"00", x"2e", x"2e", x"2e", x"32", x"2e", x"32", x"32", x"2e", x"2e", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"04", x"04", x"04", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"29", x"2d", x"5b", x"32", x"52", x"32", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"2e", x"00", x"00", x"00", x"00", x"2e", x"2e", x"32", x"32", x"2e", x"32", x"32", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"2e", x"2e", x"32", x"00", x"00", x"00", x"00", x"2e", x"2e", x"2e", x"2e", x"2e", x"2e", x"2d", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"32", x"32", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"52", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"09", x"09", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"29", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"09", x"09", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"2d", x"09", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"2e", x"2d", x"2d", x"2e", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"09", x"2e", x"32", x"32", x"2e", x"09", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"09", x"56", x"5b", x"5b", x"5b", x"5b", x"56", x"05", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"09", x"09", x"09", x"04", x"00", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"29", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"04", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"32", x"32", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"04", x"32", x"56", x"5b", x"5b", x"56", x"32", x"04", x"00", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"05", x"09", x"09", x"09", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"29", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"32", x"32", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"2e", x"2d", x"2d", x"2e", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2e", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"00", x"2d", x"00", x"00", x"00", x"2e", x"09", x"00", x"00", x"00", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"32", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"32", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"29", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"05", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"2d", x"00", x"00", x"00", x"00", x"5b", x"5b", x"04", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"32", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"2e", x"2d", x"2d", x"2d", x"2e", x"56", x"5b", x"5b", x"5b", x"5b", x"32", x"56", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2d", x"5b", x"5b", x"5b", x"00", x"00", x"04", x"56", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"56", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2e", x"5b", x"2e", x"00", x"00", x"00", x"2e", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"32", x"00", x"00", x"00", x"09", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"2d", x"32", x"32", x"32", x"2d", x"00", x"00", x"00", x"00", x"5b", x"5b", x"00", x"00", x"00", x"00", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"00", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"04", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"29", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"00", x"00", x"52", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"09", x"00", x"00", x"29", x"32", x"32", x"32", x"2d", x"00", x"00", x"09", x"32", x"32", x"2e", x"04", x"00", x"00", x"00", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2d", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"32", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"56", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"2d", x"32", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"04", x"04", x"04", x"5b", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"56", x"56", x"5b", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2d", x"2d", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"52", x"00", x"00", x"09", x"56", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"56", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"09", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"32", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"2e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"29", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"32", x"2d", x"29", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"), 
	(x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b", x"5b"));
	
	
end local_display;
